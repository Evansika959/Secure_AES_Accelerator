typedef enum logic [1:0] {
    INVALID,
    ENCRYPT,
    DECRYPT
} job_t;