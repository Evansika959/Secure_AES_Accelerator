/afs/umich.edu/class/eecs627/ibm13/artisan/2005q3v1/aci/sc-x/lef/ibm13rvt_macros.lef